-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 64-Bit"
-- VERSION		"Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"
-- CREATED		"Sun Mar 28 10:11:09 2021"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Add32 IS 
	PORT
	(
		R1 :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		R2 :  IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
		OVERFLOW :  OUT  STD_LOGIC;
		RES :  OUT  STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END Add32;

ARCHITECTURE bdf_type OF Add32 IS 

COMPONENT add
	PORT(CARRY : IN STD_LOGIC;
		 R1 : IN STD_LOGIC;
		 R2 : IN STD_LOGIC;
		 OVERFLOW : OUT STD_LOGIC;
		 RESULT : OUT STD_LOGIC
	);
END COMPONENT;

SIGNAL	RES_ALTERA_SYNTHESIZED :  STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_5 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_24 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_25 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_27 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_28 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_29 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_30 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_31 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_0 <= '0';



b2v_add0 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_0,
		 R1 => R1(0),
		 R2 => R2(0),
		 OVERFLOW => SYNTHESIZED_WIRE_1,
		 RESULT => RES_ALTERA_SYNTHESIZED(0));


b2v_add1 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_1,
		 R1 => R1(1),
		 R2 => R2(1),
		 OVERFLOW => SYNTHESIZED_WIRE_12,
		 RESULT => RES_ALTERA_SYNTHESIZED(1));


b2v_add10 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_2,
		 R1 => R1(10),
		 R2 => R2(10),
		 OVERFLOW => SYNTHESIZED_WIRE_3,
		 RESULT => RES_ALTERA_SYNTHESIZED(10));


b2v_add11 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_3,
		 R1 => R1(11),
		 R2 => R2(11),
		 OVERFLOW => SYNTHESIZED_WIRE_4,
		 RESULT => RES_ALTERA_SYNTHESIZED(11));


b2v_add12 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_4,
		 R1 => R1(12),
		 R2 => R2(12),
		 OVERFLOW => SYNTHESIZED_WIRE_5,
		 RESULT => RES_ALTERA_SYNTHESIZED(12));


b2v_add13 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_5,
		 R1 => R1(13),
		 R2 => R2(13),
		 OVERFLOW => SYNTHESIZED_WIRE_6,
		 RESULT => RES_ALTERA_SYNTHESIZED(13));


b2v_add14 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_6,
		 R1 => R1(14),
		 R2 => R2(14),
		 OVERFLOW => SYNTHESIZED_WIRE_7,
		 RESULT => RES_ALTERA_SYNTHESIZED(14));


b2v_add15 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_7,
		 R1 => R1(15),
		 R2 => R2(15),
		 OVERFLOW => SYNTHESIZED_WIRE_8,
		 RESULT => RES_ALTERA_SYNTHESIZED(15));


b2v_add16 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_8,
		 R1 => R1(16),
		 R2 => R2(16),
		 OVERFLOW => SYNTHESIZED_WIRE_9,
		 RESULT => RES_ALTERA_SYNTHESIZED(16));


b2v_add17 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_9,
		 R1 => R1(17),
		 R2 => R2(17),
		 OVERFLOW => SYNTHESIZED_WIRE_10,
		 RESULT => RES_ALTERA_SYNTHESIZED(17));


b2v_add18 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_10,
		 R1 => R1(18),
		 R2 => R2(18),
		 OVERFLOW => SYNTHESIZED_WIRE_11,
		 RESULT => RES_ALTERA_SYNTHESIZED(18));


b2v_add19 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_11,
		 R1 => R1(19),
		 R2 => R2(19),
		 OVERFLOW => SYNTHESIZED_WIRE_13,
		 RESULT => RES_ALTERA_SYNTHESIZED(19));


b2v_add2 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_12,
		 R1 => R1(2),
		 R2 => R2(2),
		 OVERFLOW => SYNTHESIZED_WIRE_23,
		 RESULT => RES_ALTERA_SYNTHESIZED(2));


b2v_add20 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_13,
		 R1 => R1(20),
		 R2 => R2(20),
		 OVERFLOW => SYNTHESIZED_WIRE_14,
		 RESULT => RES_ALTERA_SYNTHESIZED(20));


b2v_add21 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_14,
		 R1 => R1(21),
		 R2 => R2(21),
		 OVERFLOW => SYNTHESIZED_WIRE_15,
		 RESULT => RES_ALTERA_SYNTHESIZED(21));


b2v_add22 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_15,
		 R1 => R1(22),
		 R2 => R2(22),
		 OVERFLOW => SYNTHESIZED_WIRE_16,
		 RESULT => RES_ALTERA_SYNTHESIZED(22));


b2v_add23 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_16,
		 R1 => R1(23),
		 R2 => R2(23),
		 OVERFLOW => SYNTHESIZED_WIRE_17,
		 RESULT => RES_ALTERA_SYNTHESIZED(23));


b2v_add24 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_17,
		 R1 => R1(24),
		 R2 => R2(24),
		 OVERFLOW => SYNTHESIZED_WIRE_18,
		 RESULT => RES_ALTERA_SYNTHESIZED(24));


b2v_add25 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_18,
		 R1 => R1(25),
		 R2 => R2(25),
		 OVERFLOW => SYNTHESIZED_WIRE_19,
		 RESULT => RES_ALTERA_SYNTHESIZED(25));


b2v_add26 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_19,
		 R1 => R1(26),
		 R2 => R2(26),
		 OVERFLOW => SYNTHESIZED_WIRE_20,
		 RESULT => RES_ALTERA_SYNTHESIZED(26));


b2v_add27 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_20,
		 R1 => R1(27),
		 R2 => R2(27),
		 OVERFLOW => SYNTHESIZED_WIRE_21,
		 RESULT => RES_ALTERA_SYNTHESIZED(27));


b2v_add28 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_21,
		 R1 => R1(28),
		 R2 => R2(28),
		 OVERFLOW => SYNTHESIZED_WIRE_22,
		 RESULT => RES_ALTERA_SYNTHESIZED(28));


b2v_add29 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_22,
		 R1 => R1(29),
		 R2 => R2(29),
		 OVERFLOW => SYNTHESIZED_WIRE_24,
		 RESULT => RES_ALTERA_SYNTHESIZED(29));


b2v_add3 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_23,
		 R1 => R1(3),
		 R2 => R2(3),
		 OVERFLOW => SYNTHESIZED_WIRE_26,
		 RESULT => RES_ALTERA_SYNTHESIZED(3));


b2v_add30 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_24,
		 R1 => R1(30),
		 R2 => R2(30),
		 OVERFLOW => SYNTHESIZED_WIRE_25,
		 RESULT => RES_ALTERA_SYNTHESIZED(30));


b2v_add31 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_25,
		 R1 => R1(31),
		 R2 => R2(31),
		 OVERFLOW => OVERFLOW,
		 RESULT => RES_ALTERA_SYNTHESIZED(31));


b2v_add4 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_26,
		 R1 => R1(4),
		 R2 => R2(4),
		 OVERFLOW => SYNTHESIZED_WIRE_27,
		 RESULT => RES_ALTERA_SYNTHESIZED(4));


b2v_add5 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_27,
		 R1 => R1(5),
		 R2 => R2(5),
		 OVERFLOW => SYNTHESIZED_WIRE_28,
		 RESULT => RES_ALTERA_SYNTHESIZED(5));


b2v_add6 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_28,
		 R1 => R1(6),
		 R2 => R2(6),
		 OVERFLOW => SYNTHESIZED_WIRE_29,
		 RESULT => RES_ALTERA_SYNTHESIZED(6));


b2v_add7 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_29,
		 R1 => R1(7),
		 R2 => R2(7),
		 OVERFLOW => SYNTHESIZED_WIRE_30,
		 RESULT => RES_ALTERA_SYNTHESIZED(7));


b2v_add8 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_30,
		 R1 => R1(8),
		 R2 => R2(8),
		 OVERFLOW => SYNTHESIZED_WIRE_31,
		 RESULT => RES_ALTERA_SYNTHESIZED(8));


b2v_add9 : add
PORT MAP(CARRY => SYNTHESIZED_WIRE_31,
		 R1 => R1(9),
		 R2 => R2(9),
		 OVERFLOW => SYNTHESIZED_WIRE_2,
		 RESULT => RES_ALTERA_SYNTHESIZED(9));


RES <= RES_ALTERA_SYNTHESIZED;

END bdf_type;